* Extracted by KLayout with GF180MCU LVS runset on : 25/09/2025 18:50

.SUBCKT TOP
M$1 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$2 VIN_INT VIN_INT \$267 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$3 \$250 VIN_INT \$249 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$4 \$252 VIN_INT \$251 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$5 \$254 VIN_INT \$253 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$6 VIN_OUT VIN_INT \$255 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$7 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$8 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$9 \$267 \$267 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$10 \$249 \$267 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$11 \$251 \$267 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$12 \$253 \$267 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$13 \$255 \$267 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$14 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$15 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$16 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$17 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$18 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$19 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$20 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$21 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$22 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$23 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$24 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$25 VBIAS_INT VBIAS_INT \$356 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P
+ PS=21.2U PD=21.2U
M$26 \$358 VBIAS_INT \$357 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$27 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$28 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$29 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$30 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$31 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$32 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$33 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$34 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$35 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$36 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$37 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$38 \$349 \$349 \$360 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$39 \$316 \$349 \$361 VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$40 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$41 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$42 \$267 ENA VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$43 \$267 ENA VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$44 \$267 ENA VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$45 \$267 ENA VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$46 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$47 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$48 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$49 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$50 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$51 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$52 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$53 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$54 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$55 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$56 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$57 \$356 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$58 \$357 \$356 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$59 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$60 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$61 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$62 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$63 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$64 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$65 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$66 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$67 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$68 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$69 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$70 \$360 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$71 \$361 \$360 VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$72 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$73 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$74 \$356 ENA VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$75 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$76 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$77 \$360 ENA VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=6P AD=6P PS=21.2U
+ PD=21.2U
M$78 VDD|VSS VDD|VSS VDD|VSS VDD|VSS pfet_03v3 L=2U W=10U AS=5.8P AD=5.8P
+ PS=21.16U PD=21.16U
M$79 VDD|VSS IE|PD \$203 \$206 pfet_05v0 L=0.5U W=0.9U AS=0.396P AD=0.396P
+ PS=2.68U PD=2.68U
M$80 VDD|VSS \$150 \$150 \$215 pfet_05v0 L=0.5U W=0.9U AS=0.396P AD=0.396P
+ PS=2.68U PD=2.68U
M$81 VDD|VSS VDD|VSS VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P
+ PS=17.16U PD=17.16U
M$82 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$83 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$84 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$85 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$86 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$87 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$88 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$89 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$90 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$91 \$359 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$92 \$370 \$359 VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$93 VDD|VSS VDD|VSS VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P
+ PS=17.16U PD=17.16U
M$94 VDD|VSS VDD|VSS VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P AD=4.64P
+ PS=17.16U PD=17.16U
M$95 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$96 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$97 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$98 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$99 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$100 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$101 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$102 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$103 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$104 \$358 \$358 \$359 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$105 \$349 \$358 \$370 gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.8P AD=4.8P
+ PS=17.2U PD=17.2U
M$106 VDD|VSS VDD|VSS VDD|VSS gf180mcu_gnd nfet_03v3 L=1U W=8U AS=4.64P
+ AD=4.64P PS=17.16U PD=17.16U
M$107 VDD|VSS IE|PD IE|PD gf180mcu_gnd nfet_05v0 L=0.6U W=0.66U AS=0.2904P
+ AD=0.2904P PS=2.2U PD=2.2U
M$108 VDD|VSS \$150 \$212 gf180mcu_gnd nfet_05v0 L=0.6U W=0.66U AS=0.2904P
+ AD=0.2904P PS=2.2U PD=2.2U
M$109 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$110 \$250 \$250 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$111 VCM_OUT \$250 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$112 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$113 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$114 \$270 \$270 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$115 \$290 \$270 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$116 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$117 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$118 \$252 \$252 \$270 VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$119 BCM_OUT \$252 \$290 VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$120 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$121 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$122 CCM_OUT \$316 \$314 VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$123 \$316 \$314 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$124 CCM_OUT \$316 \$314 VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$125 \$316 \$314 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$126 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$127 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$128 \$350 \$254 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$129 \$314 \$254 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$130 \$350 \$254 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$131 \$314 \$254 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$132 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$133 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
M$134 \$316 \$350 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$135 \$254 \$316 \$350 VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$136 \$316 \$350 VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P
+ PS=9.2U PD=9.2U
M$137 \$254 \$316 \$350 VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.4P AD=2.4P PS=9.2U
+ PD=9.2U
M$138 VDD|VSS VDD|VSS VDD|VSS VDD|VSS nfet_03v3_dn L=1U W=4U AS=2.32P AD=2.32P
+ PS=9.16U PD=9.16U
D$139 VDD|VSS ENA diode_nd2ps_06v0 A=100P P=40U
D$140 VDD|VSS ENA diode_nd2ps_06v0 A=100P P=40U
D$141 VDD|VSS ENA diode_nd2ps_06v0 A=100P P=40U
D$142 VDD|VSS ENA diode_nd2ps_06v0 A=100P P=40U
D$143 VDD|VSS VBIAS_INT diode_nd2ps_06v0 A=100P P=40U
D$144 VDD|VSS VBIAS_INT diode_nd2ps_06v0 A=100P P=40U
D$145 VDD|VSS VBIAS_INT diode_nd2ps_06v0 A=100P P=40U
D$146 VDD|VSS VBIAS_INT diode_nd2ps_06v0 A=100P P=40U
D$147 VDD|VSS VIN_INT diode_nd2ps_06v0 A=100P P=40U
D$148 VDD|VSS VIN_INT diode_nd2ps_06v0 A=100P P=40U
D$149 VDD|VSS VIN_INT diode_nd2ps_06v0 A=100P P=40U
D$150 VDD|VSS VIN_INT diode_nd2ps_06v0 A=100P P=40U
D$151 ENA VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$152 ENA VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$153 ENA VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$154 ENA VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$155 VBIAS_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$156 VBIAS_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$157 VBIAS_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$158 VBIAS_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$159 VIN_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$160 VIN_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$161 VIN_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
D$162 VIN_INT VDD|VSS diode_pd2nw_06v0 A=100P P=40U
R$163 ENA EN gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
R$164 VBIAS_INT VBIAS gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
R$165 VIN_INT VIN gf180mcu_gnd 87.5 ppolyf_u L=10U W=40U
.ENDS TOP
